// ==================================================
//	[ VLSISYS Lab. ]
//	* Author		: Woong Choi (woongchoi@sm.ac.kr)
//	* Filename		: temp.v
//	* Description	: 
// ==================================================


module module_name(o_data, o_valid, i_data, i_ctrl);
	output reg	[BW_DATA-1:0]	o_data  ;
	output reg					o_valid ;
	input		[BW_DATA-1:0]	i_data  ;
	input		[BW_CTRL-1:0]	i_ctrl  ;

	// description of module

endmodule

module module_name
(	
	output reg	[BW_DATA-1:0]	o_data,
	output reg					o_valid,
	input		[BW_DATA-1:0]	i_data,
	input		[BW_CTRL-1:0]	i_ctrl
);

	// description of module

endmodule

